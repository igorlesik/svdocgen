import MyPkg::*;

class MyClass;
    ETrafficLight light;
endclass